* Created by KLayout

* cell a
.SUBCKT a
* net 16 vdda
* net 17 inp
* net 19 inn
* net 21 vssa
* device instance $1 r0 *1 121.5,307.5 NMOS
M$1 21 3 4 21 NMOS L=1U W=5U AS=10P AD=10P PS=14U PD=14U
* device instance $2 r0 *1 121.5,322.5 PMOS
M$2 16 3 4 16 PMOS L=1U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $3 r0 *1 14.6,348 NMOS
M$3 6 14 14 21 NMOS L=1.2U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $4 m90 *1 7.4,348 NMOS
M$4 8 14 11 21 NMOS L=1.2U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $5 m0 *1 15.6,387 PMOS
M$5 14 11 16 16 PMOS L=1.2U W=108U AS=162P AD=162P PS=168U PD=168U
* device instance $7 r180 *1 6.4,387 PMOS
M$7 11 11 16 16 PMOS L=1.2U W=108U AS=162P AD=162P PS=168U PD=168U
* device instance $9 m90 *1 110.4,317 NMOS
M$9 21 3 1 21 NMOS L=1.2U W=24U AS=48P AD=48P PS=52U PD=52U
* device instance $10 m90 *1 7.4,319 NMOS
M$10 1 6 8 21 NMOS L=1.2U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $11 r0 *1 14.6,319 NMOS
M$11 21 6 6 21 NMOS L=1.2U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $12 r0 *1 72.1,399 PMOS
M$12 16 18 9 16 PMOS L=1.2U W=36U AS=72P AD=72P PS=76U PD=76U
* device instance $13 m90 *1 62.9,399 PMOS
M$13 16 18 18 16 PMOS L=1.2U W=36U AS=72P AD=72P PS=76U PD=76U
* device instance $14 r0 *1 44.1,331 NMOS
M$14 21 12 13 21 NMOS L=1.2U W=54U AS=108P AD=108P PS=112U PD=112U
* device instance $15 m90 *1 29.9,331 NMOS
M$15 21 12 12 21 NMOS L=1.2U W=54U AS=108P AD=108P PS=112U PD=112U
* device instance $16 r0 *1 37.1,331 NMOS
M$16 21 12 15 21 NMOS L=1.2U W=54U AS=108P AD=108P PS=112U PD=112U
* device instance $17 r180 *1 126.6,394 PMOS
M$17 10 2 16 16 PMOS L=1.2U W=240U AS=280P AD=280P PS=294U PD=294U
* device instance $23 m0 *1 83.7,394 PMOS
M$23 5 9 16 16 PMOS L=1.2U W=240U AS=280P AD=280P PS=294U PD=294U
* device instance $29 m0 *1 135.6,329.5 NMOS
M$29 10 2 21 21 NMOS L=1.2U W=180U AS=225P AD=225P PS=235U PD=235U
* device instance $33 r0 *1 91.1,336.6 NMOS
M$33 21 12 5 21 NMOS L=1.2U W=180U AS=225P AD=225P PS=235U PD=235U
* device instance $37 r90 *1 117,359.5 PMOS
M$37 5 4 2 16 PMOS L=1U W=20U AS=30P AD=30P PS=36U PD=36U
* device instance $39 m0 *1 29.6,400.5 PMOS
M$39 12 11 16 16 PMOS L=1.2U W=54U AS=81P AD=81P PS=87U PD=87U
* device instance $41 r0 *1 42.1,382 PMOS
M$41 20 15 15 16 PMOS L=1.2U W=72U AS=90P AD=90P PS=100U PD=100U
* device instance $45 r0 *1 42.1,408 PMOS
M$45 16 20 20 16 PMOS L=1.2U W=72U AS=90P AD=90P PS=100U PD=100U
* device instance $49 m90 *1 71.4,369 NMOS
M$49 13 19 9 21 NMOS L=1.2U W=6U AS=12P AD=12P PS=16U PD=16U
* device instance $50 r0 *1 64.1,369 NMOS
M$50 13 17 18 21 NMOS L=1.2U W=6U AS=12P AD=12P PS=16U PD=16U
* device instance $51 r270 *1 64.3,321.6 CAP
C$51 7 5 1.032e-012
* device instance $52 r270 *1 145,397.7 CAP
C$52 5 10 1.032e-012
* device instance $53 m45 *1 68.65,347.4 PMOS
M$53 7 15 9 16 PMOS L=1.2U W=55U AS=82.5P AD=82.5P PS=88.5U PD=88.5U
* device instance $55 r180 *1 123.5,341.5 NMOS
M$55 2 4 21 21 NMOS L=1U W=12U AS=18P AD=18P PS=24U PD=24U
* device instance $57 r90 *1 118,351 NMOS
M$57 2 3 5 21 NMOS L=1U W=12U AS=24P AD=24P PS=28U PD=28U
.ENDS a
