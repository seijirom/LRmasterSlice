* Z:\HOME\SEIJIROM\DROPBOX\WORK\LRMASTERSLICE\Ã‚³ÃƑ³ÃƑ‘ÃƑ¬ÃƑ¼Ã‚¿\COMP_NLF.ASC
*
.SUBCKT COMP_NLF INP INN XSTBY OUT VDDA VSSA
M6 STBY XSTBY VSSA VSSA NCH L=1.0U W=5.0U M=1
M9 VDDA XSTBY STBY VDDA PCH L=1.0U W=10.0U M=1
M_18 N001 N004 N012 VSSA NCH L=1.2U W=10.0U M=1
M_14 VDDA N001 N004 VDDA PCH L=1.2U W=108.0U M=2
M_17 VDDA N001 N001 VDDA PCH L=1.2U W=108.0U M=2
M_15 N004 N004 N011 VSSA NCH L=1.2U W=10.0U M=1
M_20 N014 XSTBY VSSA VSSA NCH L=1.2U W=24.0U M=1
M_19 N012 N011 N014 VSSA NCH L=1.2U W=30.0U M=1
M_16 N011 N011 VSSA VSSA NCH L=1.2U W=30.0U M=1
M_4 VDDA N003 N005 VDDA PCH L=1.2U W=36.0U M=1
M_5 N013 N010 VSSA VSSA NCH L=1.2U W=54.0U M=1
M_8 VDDA N005 N008 VDDA PCH L=1.2U W=240.0U M=6
M_7 N008 N010 VSSA VSSA NCH L=1.2U W=180.00U M=2
M_100 OUT N009 VSSA VSSA NCH L=1.2U W=180.0U M=2
M_101 VDDA N009 OUT VDDA PCH L=1.2U W=240.0U M=6
C2 N008 N007 1.032P
C7 OUT N008 1.032P
M29 N008 STBY N009 VDDA PCH L=1.0U W=20.0U M=1
M30 N009 XSTBY N008 VSSA NCH L=1.0U W=12.0U M=1
M31 N009 STBY VSSA VSSA NCH L=1.0U W=12.0U M=1
M_13 VDDA N001 N010 VDDA PCH L=1.2U W=54.0U M=1
M_11 VDDA N002 N002 VDDA PCH L=1.2U W=72.0U M=1
M_10 N002 N006 N006 VDDA PCH L=1.2U W=72.0U M=1
M_12 N010 N010 VSSA VSSA NCH L=1.2U W=54.0U M=1
M_9 N006 N010 VSSA VSSA NCH L=1.2U W=54.0U M=1
M_1 N003 INP N013 VSSA NCH L=1.2U W=6.0U M=1
M_2 N005 INN N013 VSSA NCH L=1.2U W=6.0U M=1
M_3 VDDA N003 N003 VDDA PCH L=1.2U W=36.0U M=1
M_6 N005 N006 N007 VDDA PCH L=1.2U W=55.0U M=1
.ENDS COMP_NLF

