* Z:\HOME\SEIJIROM\DROPBOX\WORK\LRMASTERSLICE\Ã‚³ÃƑ³ÃƑ‘ÃƑ¬ÃƑ¼Ã‚¿\COMP_PLF.ASC
*
.SUBCKT COMP_PLF INP INN XSTBY OUT VDDA VSSA
M33 VBP_B VBN_B N007 VSSA NCH L=1.2U W=6.45U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M34 NC_01 VBP_B VBN_B VDDA PCH L=1.2U W=13.8U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M37 VDDA VBP_B VBP_B VDDA PCH L=1.2U W=13.8U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M38 VBN_B VBN_B N006 VSSA NCH L=1.2U W=6.45U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M39 N010 XSTBY VSSA VSSA NCH L=2.0U W=3.3U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M40 N007 N006 N010 VSSA NCH L=1.2U W=18.1U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M41 N006 N006 VSSA VSSA NCH L=1.2U W=7.2U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M42 VDDA VBP_B N001 VDDA PCH L=1.2U W=13.5U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M43 N008 N009 VSSA VSSA NCH L=1.2U W=3.7U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M44 N009 N009 VSSA VSSA NCH L=1.2U W=3.7U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M45 N001 INN N008 N001 PCH L=1.2U W=10.0U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M46 N001 INP N009 N001 PCH L=1.2U W=10.0U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M47 VDDA VBP_B N003 VDDA PCH L=1.2U W=200.0U PD=W+L+L PS=PD AD=W*L AS=AD M=10
M48 N003 N008 VSSA VSSA NCH L=1.2U W=95.2U PD=W+L+L PS=PD AD=W*L AS=AD M=4
M49 OUT N005 VSSA VSSA NCH L=1.2U W=24.66U PD=W+L+L PS=PD AD=W*L AS=AD M=2
M50 VDDA N005 OUT VDDA PCH L=1.2U W=80.0U PD=W+L+L PS=PD AD=W*L AS=AD M=4
C4 N003 N002 1P
C5 OUT VSSA 1P
C6 OUT N003 1P
M1 N003 N004 N005 VDDA PCH L=1.0U W=20.0U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M2 N005 XSTBY N003 VSSA NCH L=1.0U W=12.0U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M3 N004 XSTBY VSSA VSSA NCH L=1.0U W=12.0U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M4 VDDA XSTBY N004 VDDA PCH L=1.0U W=20.0U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M5 N005 N004 VSSA VSSA NCH L=1.0U W=12.0U PD=W+L+L PS=PD AD=W*L AS=AD M=1
M6 N008 VBN_B N002 VSSA NCH L=1.2U W=28.8U PD=W+L+L PS=PD AD=W*L AS=AD M=2
.ENDS COMP_PLF

