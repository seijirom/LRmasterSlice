* C:\USERS\SEIJIROM\DROPBOX\WORK\LRMASTERSLICE\³0Ó0Ñ0Ì0Ü0¿0\COMP_NLF.ASC
*
.SUBCKT COMP_NLF INP INN XSTBY OUT VDDA VSSA
M6 STBY XSTBY VSSA VSSA NCH L=1.0U W=5.0U M=1
M9 VDDA XSTBY STBY VDDA PCH L=1.0U W=10.0U M=1
M_18 N002 N005 N014 VSSA NCH L=1.2U W=10.0U M=1
M_14 N001 N002 N005 N001 PCH L=1.2U W=108.0U M=2
M_17 N001 N002 N002 N001 PCH L=1.2U W=108.0U M=2
M_15 N005 N005 N013 VSSA NCH L=1.2U W=10.0U M=1
M_20 N016 XSTBY VSSA VSSA NCH L=1.2U W=24.0U M=1
M_19 N014 N013 N016 VSSA NCH L=1.2U W=30.0U M=1
M_16 N013 N013 VSSA VSSA NCH L=1.2U W=30.0U M=1
M_4 N001 N004 N006 N001 PCH L=1.2U W=36.0U M=1
M_5 N015 N012 VSSA VSSA NCH L=1.2U W=54.0U M=1
M_8 N001 N006 N009 N001 PCH L=1.2U W=240.0U M=6
M_7 N009 N012 VSSA VSSA NCH L=1.2U W=180.16U M=2
M_100 OUT N011 VSSA VSSA NCH L=1.2U W=180.0U M=2
M_101 N001 N011 OUT N001 PCH L=1.2U W=240.0U M=6
C2 N009 N008 1P
C7 OUT N009 1P
M29 N009 STBY N011 N001 PCH L=1.0U W=20.0U M=1
M30 N011 XSTBY N009 VSSA NCH L=1.0U W=12.0U M=1
M31 N011 STBY VSSA VSSA NCH L=1.0U W=12.0U M=1
M_13 N001 N002 N012 N001 PCH L=1.2U W=54.0U M=1
M_11 N001 N003 N003 N001 PCH L=1.2U W=72.0U M=1
M_10 N003 N007 N007 N001 PCH L=1.2U W=72.0U M=1
M_12 N012 N012 VSSA VSSA NCH L=1.2U W=54.0U M=1
M_9 N007 N012 VSSA VSSA NCH L=1.2U W=54.0U M=1
M_1 N004 INP N015 N010 NCH L=1.2U W=6.0U M=1
M_2 N006 INN N015 N010 NCH L=1.2U W=6.0U M=1
M_3 N001 N004 N004 N001 PCH L=1.2U W=36.0U M=1
M_6 N006 N007 N008 N001 PCH L=1.2U W=55.0U M=1
R2 N001 VDDA 0.01
.ENDS COMP_NLF

